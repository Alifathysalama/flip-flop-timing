magic
tech ihp-sg13g2
timestamp 1758009537
<< nwell >>
rect -69 0 1100 148
<< nmos >>
rect 0 -61 13 -31
rect 31 -61 44 -31
rect 82 -61 95 -31
rect 214 -61 227 -31
rect 245 -61 258 -31
rect 370 -61 383 -31
rect 410 -61 423 -31
rect 449 -61 462 -31
rect 574 -61 587 -31
rect 615 -61 628 -31
rect 656 -61 669 -31
rect 762 -61 775 -31
rect 801 -61 814 -31
rect 841 -61 854 -31
rect 966 -61 979 -31
rect 997 -61 1010 -31
<< pmos >>
rect 0 31 13 61
rect 51 31 64 61
rect 102 31 115 61
rect 204 31 217 61
rect 255 31 268 61
rect 347 31 360 61
rect 398 31 411 61
rect 449 31 462 61
rect 551 31 564 61
rect 602 31 615 61
rect 653 31 666 61
rect 762 31 775 61
rect 813 31 826 61
rect 864 31 877 61
rect 966 31 979 61
rect 1017 31 1030 61
<< ndiff >>
rect -34 -38 0 -31
rect -34 -54 -27 -38
rect -11 -54 0 -38
rect -34 -61 0 -54
rect 13 -61 31 -31
rect 44 -61 82 -31
rect 95 -38 129 -31
rect 95 -54 106 -38
rect 122 -54 129 -38
rect 95 -61 129 -54
rect 180 -38 214 -31
rect 180 -54 187 -38
rect 203 -54 214 -38
rect 180 -61 214 -54
rect 227 -61 245 -31
rect 258 -38 292 -31
rect 258 -54 269 -38
rect 285 -54 292 -38
rect 258 -61 292 -54
rect 336 -38 370 -31
rect 336 -54 343 -38
rect 359 -54 370 -38
rect 336 -61 370 -54
rect 383 -61 410 -31
rect 423 -61 449 -31
rect 462 -38 496 -31
rect 462 -54 473 -38
rect 489 -54 496 -38
rect 462 -61 496 -54
rect 540 -38 574 -31
rect 540 -54 547 -38
rect 563 -54 574 -38
rect 540 -61 574 -54
rect 587 -61 615 -31
rect 628 -61 656 -31
rect 669 -38 703 -31
rect 669 -54 680 -38
rect 696 -54 703 -38
rect 669 -61 703 -54
rect 728 -38 762 -31
rect 728 -54 735 -38
rect 751 -54 762 -38
rect 728 -61 762 -54
rect 775 -61 801 -31
rect 814 -61 841 -31
rect 854 -38 888 -31
rect 854 -54 865 -38
rect 881 -54 888 -38
rect 854 -61 888 -54
rect 932 -38 966 -31
rect 932 -54 939 -38
rect 955 -54 966 -38
rect 932 -61 966 -54
rect 979 -61 997 -31
rect 1010 -38 1044 -31
rect 1010 -54 1021 -38
rect 1037 -54 1044 -38
rect 1010 -61 1044 -54
<< pdiff >>
rect -34 54 0 61
rect -34 38 -27 54
rect -11 38 0 54
rect -34 31 0 38
rect 13 54 51 61
rect 13 38 24 54
rect 40 38 51 54
rect 13 31 51 38
rect 64 54 102 61
rect 64 38 75 54
rect 91 38 102 54
rect 64 31 102 38
rect 115 54 149 61
rect 115 38 126 54
rect 142 38 149 54
rect 115 31 149 38
rect 170 54 204 61
rect 170 38 177 54
rect 193 38 204 54
rect 170 31 204 38
rect 217 54 255 61
rect 217 38 228 54
rect 244 38 255 54
rect 217 31 255 38
rect 268 54 347 61
rect 268 38 279 54
rect 295 38 320 54
rect 336 38 347 54
rect 268 31 347 38
rect 360 54 398 61
rect 360 38 371 54
rect 387 38 398 54
rect 360 31 398 38
rect 411 54 449 61
rect 411 38 422 54
rect 438 38 449 54
rect 411 31 449 38
rect 462 54 496 61
rect 462 38 473 54
rect 489 38 496 54
rect 462 31 496 38
rect 517 54 551 61
rect 517 38 524 54
rect 540 38 551 54
rect 517 31 551 38
rect 564 54 602 61
rect 564 38 575 54
rect 591 38 602 54
rect 564 31 602 38
rect 615 54 653 61
rect 615 38 626 54
rect 642 38 653 54
rect 615 31 653 38
rect 666 54 701 61
rect 666 38 677 54
rect 693 38 701 54
rect 666 31 701 38
rect 728 54 762 61
rect 728 38 735 54
rect 751 38 762 54
rect 728 31 762 38
rect 775 54 813 61
rect 775 38 786 54
rect 802 38 813 54
rect 775 31 813 38
rect 826 54 864 61
rect 826 38 837 54
rect 853 38 864 54
rect 826 31 864 38
rect 877 54 911 61
rect 877 38 888 54
rect 904 38 911 54
rect 877 31 911 38
rect 932 54 966 61
rect 932 38 939 54
rect 955 38 966 54
rect 932 31 966 38
rect 979 54 1017 61
rect 979 38 990 54
rect 1006 38 1017 54
rect 979 31 1017 38
rect 1030 54 1065 61
rect 1030 38 1041 54
rect 1057 38 1065 54
rect 1030 31 1065 38
<< ndiffc >>
rect -27 -54 -11 -38
rect 106 -54 122 -38
rect 187 -54 203 -38
rect 269 -54 285 -38
rect 343 -54 359 -38
rect 473 -54 489 -38
rect 547 -54 563 -38
rect 680 -54 696 -38
rect 735 -54 751 -38
rect 865 -54 881 -38
rect 939 -54 955 -38
rect 1021 -54 1037 -38
<< pdiffc >>
rect -27 38 -11 54
rect 24 38 40 54
rect 75 38 91 54
rect 126 38 142 54
rect 177 38 193 54
rect 228 38 244 54
rect 279 38 295 54
rect 320 38 336 54
rect 371 38 387 54
rect 422 38 438 54
rect 473 38 489 54
rect 524 38 540 54
rect 575 38 591 54
rect 626 38 642 54
rect 677 38 693 54
rect 735 38 751 54
rect 786 38 802 54
rect 837 38 853 54
rect 888 38 904 54
rect 939 38 955 54
rect 990 38 1006 54
rect 1041 38 1057 54
<< psubdiff >>
rect -45 -101 1076 -94
rect -45 -117 -38 -101
rect -22 -117 -2 -101
rect 14 -117 34 -101
rect 51 -117 70 -101
rect 87 -117 106 -101
rect 123 -117 142 -101
rect 159 -117 178 -101
rect 195 -117 214 -101
rect 231 -117 250 -101
rect 267 -117 286 -101
rect 303 -117 322 -101
rect 339 -117 358 -101
rect 375 -117 394 -101
rect 411 -117 430 -101
rect 447 -117 466 -101
rect 483 -117 502 -101
rect 519 -117 538 -101
rect 555 -117 574 -101
rect 591 -117 610 -101
rect 627 -117 646 -101
rect 663 -117 682 -101
rect 699 -117 718 -101
rect 735 -117 754 -101
rect 771 -117 790 -101
rect 807 -117 826 -101
rect 843 -117 862 -101
rect 879 -117 898 -101
rect 915 -117 934 -101
rect 951 -117 970 -101
rect 987 -117 1006 -101
rect 1023 -117 1042 -101
rect 1059 -117 1076 -101
rect -45 -124 1076 -117
<< nsubdiff >>
rect -45 117 1076 124
rect -45 101 -38 117
rect -22 101 -2 117
rect 14 101 34 117
rect 51 101 70 117
rect 86 101 106 117
rect 122 101 142 117
rect 158 101 178 117
rect 194 101 214 117
rect 230 101 250 117
rect 266 101 286 117
rect 302 101 322 117
rect 338 101 358 117
rect 374 101 394 117
rect 410 101 430 117
rect 446 101 466 117
rect 482 101 502 117
rect 518 101 538 117
rect 554 101 574 117
rect 590 101 610 117
rect 626 101 646 117
rect 662 101 682 117
rect 698 101 718 117
rect 734 101 754 117
rect 770 101 790 117
rect 806 101 826 117
rect 842 101 862 117
rect 878 101 898 117
rect 914 101 934 117
rect 950 101 970 117
rect 986 101 1006 117
rect 1022 101 1042 117
rect 1058 101 1076 117
rect -45 94 1076 101
<< psubdiffcont >>
rect -38 -117 -22 -101
rect -2 -117 14 -101
rect 34 -117 51 -101
rect 70 -117 87 -101
rect 106 -117 123 -101
rect 142 -117 159 -101
rect 178 -117 195 -101
rect 214 -117 231 -101
rect 250 -117 267 -101
rect 286 -117 303 -101
rect 322 -117 339 -101
rect 358 -117 375 -101
rect 394 -117 411 -101
rect 430 -117 447 -101
rect 466 -117 483 -101
rect 502 -117 519 -101
rect 538 -117 555 -101
rect 574 -117 591 -101
rect 610 -117 627 -101
rect 646 -117 663 -101
rect 682 -117 699 -101
rect 718 -117 735 -101
rect 754 -117 771 -101
rect 790 -117 807 -101
rect 826 -117 843 -101
rect 862 -117 879 -101
rect 898 -117 915 -101
rect 934 -117 951 -101
rect 970 -117 987 -101
rect 1006 -117 1023 -101
rect 1042 -117 1059 -101
<< nsubdiffcont >>
rect -38 101 -22 117
rect -2 101 14 117
rect 34 101 51 117
rect 70 101 86 117
rect 106 101 122 117
rect 142 101 158 117
rect 178 101 194 117
rect 214 101 230 117
rect 250 101 266 117
rect 286 101 302 117
rect 322 101 338 117
rect 358 101 374 117
rect 394 101 410 117
rect 430 101 446 117
rect 466 101 482 117
rect 502 101 518 117
rect 538 101 554 117
rect 574 101 590 117
rect 610 101 626 117
rect 646 101 662 117
rect 682 101 698 117
rect 718 101 734 117
rect 754 101 770 117
rect 790 101 806 117
rect 826 101 842 117
rect 862 101 878 117
rect 898 101 914 117
rect 934 101 950 117
rect 970 101 986 117
rect 1006 101 1022 117
rect 1042 101 1058 117
<< poly >>
rect 0 61 13 79
rect 51 61 64 79
rect 102 61 115 79
rect 204 61 217 79
rect 255 61 268 79
rect 347 61 360 80
rect 398 61 411 80
rect 449 61 462 80
rect 551 61 564 79
rect 602 61 615 79
rect 653 61 666 79
rect 762 61 775 79
rect 813 61 826 79
rect 864 61 877 79
rect 966 61 979 79
rect 1017 61 1030 79
rect 0 15 13 31
rect 51 15 64 31
rect -21 8 13 15
rect -21 -8 -14 8
rect 2 -8 13 8
rect 34 8 64 15
rect 34 -2 41 8
rect -21 -15 13 -8
rect 0 -31 13 -15
rect 31 -8 41 -2
rect 57 -8 64 8
rect 102 17 115 31
rect 102 10 137 17
rect 102 0 114 10
rect 31 -15 64 -8
rect 100 -6 114 0
rect 130 -6 137 10
rect 100 -11 137 -6
rect 204 -11 217 31
rect 255 -11 268 31
rect 347 20 360 31
rect 330 10 360 20
rect 398 24 411 31
rect 398 14 431 24
rect 398 13 408 14
rect 330 -6 337 10
rect 353 -6 360 10
rect 330 -11 360 -6
rect 401 -2 408 13
rect 424 -2 431 14
rect 401 -9 431 -2
rect 449 15 462 31
rect 449 8 479 15
rect 449 -8 456 8
rect 472 -8 479 8
rect 82 -13 137 -11
rect 31 -31 44 -15
rect 82 -24 113 -13
rect 160 -24 227 -11
rect 82 -31 95 -24
rect 160 -31 173 -24
rect 214 -31 227 -24
rect 245 -24 312 -11
rect 330 -13 383 -11
rect 347 -24 383 -13
rect 245 -31 258 -24
rect 299 -31 312 -24
rect 370 -31 383 -24
rect 410 -31 423 -9
rect 449 -15 479 -8
rect 551 -11 564 31
rect 602 15 615 31
rect 602 8 635 15
rect 602 6 612 8
rect 605 -8 612 6
rect 628 -8 635 8
rect 449 -31 462 -15
rect 520 -24 587 -11
rect 605 -15 635 -8
rect 653 6 666 31
rect 762 15 775 31
rect 813 15 826 31
rect 864 24 877 31
rect 966 24 979 31
rect 745 8 775 15
rect 653 -1 683 6
rect 520 -31 533 -24
rect 574 -31 587 -24
rect 615 -31 628 -15
rect 653 -17 660 -1
rect 676 -17 683 -1
rect 745 -8 752 8
rect 768 -8 775 8
rect 745 -15 775 -8
rect 793 8 826 15
rect 793 -8 800 8
rect 816 6 826 8
rect 844 11 877 24
rect 926 17 979 24
rect 816 -8 823 6
rect 793 -15 823 -8
rect 844 -11 857 11
rect 926 1 933 17
rect 949 11 979 17
rect 1017 15 1030 31
rect 949 1 956 11
rect 926 -6 956 1
rect 943 -11 956 -6
rect 997 8 1035 15
rect 997 -8 1012 8
rect 1028 -8 1035 8
rect 844 -12 908 -11
rect 653 -24 683 -17
rect 656 -31 669 -24
rect 762 -31 775 -15
rect 801 -31 814 -15
rect 841 -24 908 -12
rect 943 -24 979 -11
rect 841 -31 854 -24
rect 895 -31 908 -24
rect 966 -31 979 -24
rect 997 -15 1035 -8
rect 997 -31 1010 -15
rect 136 -38 173 -31
rect 136 -54 143 -38
rect 159 -54 173 -38
rect 136 -61 173 -54
rect 299 -38 329 -31
rect 299 -54 306 -38
rect 322 -54 329 -38
rect 299 -61 329 -54
rect 503 -38 533 -31
rect 503 -54 510 -38
rect 526 -54 533 -38
rect 503 -61 533 -54
rect 895 -38 925 -31
rect 895 -54 902 -38
rect 918 -54 925 -38
rect 895 -61 925 -54
rect 0 -79 13 -61
rect 31 -79 44 -61
rect 82 -79 95 -61
rect 214 -79 227 -61
rect 245 -79 258 -61
rect 370 -79 383 -61
rect 410 -79 423 -61
rect 449 -79 462 -61
rect 574 -79 587 -61
rect 615 -79 628 -61
rect 656 -79 669 -61
rect 762 -79 775 -61
rect 801 -79 814 -61
rect 841 -79 854 -61
rect 966 -79 979 -61
rect 997 -79 1010 -61
<< polycont >>
rect -14 -8 2 8
rect 41 -8 57 8
rect 114 -6 130 10
rect 337 -6 353 10
rect 408 -2 424 14
rect 456 -8 472 8
rect 612 -8 628 8
rect 660 -17 676 -1
rect 752 -8 768 8
rect 800 -8 816 8
rect 933 1 949 17
rect 1012 -8 1028 8
rect 143 -54 159 -38
rect 306 -54 322 -38
rect 510 -54 526 -38
rect 902 -54 918 -38
<< metal1 >>
rect -45 117 1076 124
rect -45 101 -38 117
rect -22 101 -2 117
rect 14 101 34 117
rect 51 101 70 117
rect 86 101 106 117
rect 122 101 142 117
rect 158 101 178 117
rect 194 101 214 117
rect 230 101 250 117
rect 266 101 286 117
rect 302 101 322 117
rect 338 101 358 117
rect 374 101 394 117
rect 410 101 430 117
rect 446 101 466 117
rect 482 101 502 117
rect 518 101 538 117
rect 554 101 574 117
rect 590 101 610 117
rect 626 101 646 117
rect 662 101 682 117
rect 698 101 718 117
rect 734 101 754 117
rect 770 101 790 117
rect 806 101 826 117
rect 842 101 862 117
rect 878 101 898 117
rect 914 101 934 117
rect 950 101 970 117
rect 986 101 1006 117
rect 1022 101 1042 117
rect 1058 101 1076 117
rect -45 77 1076 101
rect -32 54 -4 77
rect -32 38 -27 54
rect -11 38 -4 54
rect -32 33 -4 38
rect 14 56 50 59
rect 14 36 22 56
rect 42 36 50 56
rect 14 33 50 36
rect 68 54 101 77
rect 68 38 75 54
rect 91 38 101 54
rect 68 33 101 38
rect 119 56 154 59
rect 119 36 124 56
rect 144 36 154 56
rect 119 33 154 36
rect 172 54 198 77
rect 172 38 177 54
rect 193 38 198 54
rect 172 33 198 38
rect 223 54 249 59
rect 223 38 228 54
rect 244 38 249 54
rect 223 15 249 38
rect 267 54 342 77
rect 267 38 279 54
rect 295 38 320 54
rect 336 38 342 54
rect 267 34 342 38
rect 360 56 397 59
rect 360 36 365 56
rect 385 54 397 56
rect 387 38 397 54
rect 385 36 397 38
rect 415 54 445 77
rect 415 38 422 54
rect 438 38 445 54
rect 415 36 445 38
rect 463 56 496 59
rect 463 36 471 56
rect 491 36 496 56
rect 360 35 397 36
rect 360 33 383 35
rect 463 31 496 36
rect 514 54 547 77
rect 514 38 524 54
rect 540 38 547 54
rect 514 33 547 38
rect 565 56 601 59
rect 565 36 573 56
rect 593 36 601 56
rect 565 33 601 36
rect 619 54 648 77
rect 619 38 626 54
rect 642 38 648 54
rect 619 33 648 38
rect 666 56 717 59
rect 666 36 675 56
rect 695 36 717 56
rect 401 16 431 17
rect 305 15 331 16
rect -24 10 6 15
rect -24 -10 -16 10
rect 4 -10 6 10
rect -24 -15 6 -10
rect 35 10 95 15
rect 35 8 71 10
rect 35 -8 41 8
rect 57 -8 71 8
rect 35 -10 71 -8
rect 91 -10 95 10
rect 35 -15 95 -10
rect 113 10 285 15
rect 113 -6 114 10
rect 130 -6 285 10
rect 305 -5 310 15
rect 330 10 360 15
rect 330 -5 337 10
rect 305 -6 337 -5
rect 353 -6 360 10
rect 401 -4 406 16
rect 426 -4 431 16
rect 570 13 591 33
rect 666 28 717 36
rect 735 54 758 77
rect 751 38 758 54
rect 735 33 758 38
rect 776 56 812 59
rect 776 36 784 56
rect 804 36 812 56
rect 776 33 812 36
rect 830 54 863 77
rect 830 38 837 54
rect 853 38 863 54
rect 830 33 863 38
rect 881 56 911 59
rect 881 36 886 56
rect 906 36 911 56
rect 701 15 717 28
rect 881 17 911 36
rect 929 54 960 77
rect 929 38 939 54
rect 955 38 960 54
rect 985 54 1011 59
rect 985 52 990 54
rect 929 35 960 38
rect 978 38 990 52
rect 1006 38 1011 54
rect 978 31 1011 38
rect 1029 54 1062 77
rect 1029 38 1041 54
rect 1057 38 1062 54
rect 1029 34 1062 38
rect 978 17 994 31
rect 881 15 933 17
rect 113 -12 285 -6
rect 113 -31 164 -30
rect 113 -33 122 -31
rect -32 -38 6 -33
rect -32 -54 -27 -38
rect -11 -54 6 -38
rect -32 -77 6 -54
rect 101 -38 122 -33
rect 101 -54 106 -38
rect 142 -38 164 -31
rect 142 -51 143 -38
rect 122 -54 143 -51
rect 159 -54 164 -38
rect 101 -59 164 -54
rect 182 -38 244 -33
rect 182 -54 187 -38
rect 203 -54 244 -38
rect 182 -77 244 -54
rect 262 -38 285 -12
rect 401 -15 431 -4
rect 449 8 591 13
rect 449 -8 456 8
rect 472 -8 591 8
rect 449 -13 591 -8
rect 609 10 635 15
rect 609 -10 610 10
rect 630 -10 635 10
rect 262 -54 269 -38
rect 262 -61 285 -54
rect 303 -31 325 -24
rect 609 -28 635 -10
rect 653 1 683 10
rect 653 -19 658 1
rect 678 -19 683 1
rect 653 -20 683 -19
rect 701 8 775 15
rect 701 -8 752 8
rect 768 -8 775 8
rect 701 -15 775 -8
rect 793 10 823 15
rect 793 -10 798 10
rect 818 -10 823 10
rect 793 -15 823 -10
rect 860 1 933 15
rect 949 1 954 17
rect 860 -4 954 1
rect 972 1 994 17
rect 1012 10 1048 13
rect 1012 8 1017 10
rect 303 -51 304 -31
rect 324 -51 325 -31
rect 303 -54 306 -51
rect 322 -54 325 -51
rect 303 -65 325 -54
rect 343 -38 448 -33
rect 359 -54 448 -38
rect -45 -79 244 -77
rect 343 -77 448 -54
rect 466 -36 526 -33
rect 466 -56 471 -36
rect 491 -38 526 -36
rect 491 -54 510 -38
rect 491 -56 526 -54
rect 466 -59 526 -56
rect 544 -38 591 -33
rect 701 -38 717 -15
rect 544 -54 547 -38
rect 563 -46 591 -38
rect 563 -54 651 -46
rect 544 -77 651 -54
rect 669 -54 680 -38
rect 696 -54 717 -38
rect 669 -59 717 -54
rect 735 -38 842 -33
rect 751 -54 842 -38
rect 735 -77 842 -54
rect 860 -38 884 -4
rect 972 -31 990 1
rect 1012 -10 1017 -8
rect 1037 -10 1048 10
rect 1012 -13 1048 -10
rect 860 -54 865 -38
rect 881 -54 884 -38
rect 860 -59 884 -54
rect 902 -36 990 -31
rect 902 -38 918 -36
rect 902 -56 918 -54
rect 938 -38 990 -36
rect 938 -54 939 -38
rect 955 -49 990 -38
rect 1009 -38 1044 -31
rect 955 -54 960 -49
rect 938 -56 960 -54
rect 902 -59 960 -56
rect 1009 -54 1021 -38
rect 1037 -54 1044 -38
rect 1009 -77 1044 -54
rect -45 -83 285 -79
rect 343 -83 1076 -77
rect -45 -101 1076 -83
rect -45 -117 -38 -101
rect -22 -117 -2 -101
rect 14 -117 34 -101
rect 51 -117 70 -101
rect 87 -117 106 -101
rect 123 -117 142 -101
rect 159 -117 178 -101
rect 195 -117 214 -101
rect 231 -117 250 -101
rect 267 -117 286 -101
rect 303 -117 322 -101
rect 339 -117 358 -101
rect 375 -117 394 -101
rect 411 -117 430 -101
rect 447 -117 466 -101
rect 483 -117 502 -101
rect 519 -117 538 -101
rect 555 -117 574 -101
rect 591 -117 610 -101
rect 627 -117 646 -101
rect 663 -117 682 -101
rect 699 -117 718 -101
rect 735 -117 754 -101
rect 771 -117 790 -101
rect 807 -117 826 -101
rect 843 -117 862 -101
rect 879 -117 898 -101
rect 915 -117 934 -101
rect 951 -117 970 -101
rect 987 -117 1006 -101
rect 1023 -117 1042 -101
rect 1059 -117 1076 -101
rect -45 -124 1076 -117
<< via1 >>
rect 22 54 42 56
rect 22 38 24 54
rect 24 38 40 54
rect 40 38 42 54
rect 22 36 42 38
rect 124 54 144 56
rect 124 38 126 54
rect 126 38 142 54
rect 142 38 144 54
rect 124 36 144 38
rect 365 54 385 56
rect 365 38 371 54
rect 371 38 385 54
rect 365 36 385 38
rect 471 54 491 56
rect 471 38 473 54
rect 473 38 489 54
rect 489 38 491 54
rect 471 36 491 38
rect 573 54 593 56
rect 573 38 575 54
rect 575 38 591 54
rect 591 38 593 54
rect 573 36 593 38
rect 675 54 695 56
rect 675 38 677 54
rect 677 38 693 54
rect 693 38 695 54
rect 675 36 695 38
rect -16 8 4 10
rect -16 -8 -14 8
rect -14 -8 2 8
rect 2 -8 4 8
rect -16 -10 4 -8
rect 71 -10 91 10
rect 310 -5 330 15
rect 406 14 426 16
rect 406 -2 408 14
rect 408 -2 424 14
rect 424 -2 426 14
rect 406 -4 426 -2
rect 784 54 804 56
rect 784 38 786 54
rect 786 38 802 54
rect 802 38 804 54
rect 784 36 804 38
rect 886 54 906 56
rect 886 38 888 54
rect 888 38 904 54
rect 904 38 906 54
rect 886 36 906 38
rect 122 -51 142 -31
rect 610 8 630 10
rect 610 -8 612 8
rect 612 -8 628 8
rect 628 -8 630 8
rect 610 -10 630 -8
rect 658 -1 678 1
rect 658 -17 660 -1
rect 660 -17 676 -1
rect 676 -17 678 -1
rect 658 -19 678 -17
rect 798 8 818 10
rect 798 -8 800 8
rect 800 -8 816 8
rect 816 -8 818 8
rect 798 -10 818 -8
rect 1017 8 1037 10
rect 304 -38 324 -31
rect 304 -51 306 -38
rect 306 -51 322 -38
rect 322 -51 324 -38
rect 471 -38 491 -36
rect 471 -54 473 -38
rect 473 -54 489 -38
rect 489 -54 491 -38
rect 471 -56 491 -54
rect 1017 -8 1028 8
rect 1028 -8 1037 8
rect 1017 -10 1037 -8
rect 918 -56 938 -36
<< metal2 >>
rect 323 97 532 103
rect -24 83 547 97
rect -24 77 343 83
rect 512 77 547 83
rect -24 15 -4 77
rect 364 56 496 62
rect 17 36 22 56
rect 42 36 124 56
rect 144 36 149 56
rect 364 36 365 56
rect 385 42 471 56
rect 25 31 149 36
rect -24 10 4 15
rect -24 -10 -16 10
rect -24 -15 4 -10
rect 25 -31 45 31
rect 219 10 310 15
rect 66 -10 71 10
rect 91 -5 310 10
rect 330 -5 335 15
rect 91 -10 239 -5
rect 365 -26 385 36
rect 491 36 496 56
rect 406 16 448 21
rect 426 -4 448 16
rect 406 -14 448 -4
rect 304 -31 385 -26
rect 25 -51 122 -31
rect 142 -51 283 -31
rect 260 -82 283 -51
rect 324 -46 385 -31
rect 471 -36 491 36
rect 527 10 547 77
rect 568 36 573 56
rect 593 36 675 56
rect 695 36 700 56
rect 779 36 784 56
rect 804 36 886 56
rect 906 36 911 56
rect 765 10 823 15
rect 527 -10 610 10
rect 630 -10 635 10
rect 658 1 678 6
rect 765 -10 770 10
rect 790 -10 798 10
rect 818 -10 823 10
rect 845 -10 1017 10
rect 1037 -10 1042 10
rect 658 -31 678 -19
rect 845 -31 865 -10
rect 304 -56 324 -51
rect 471 -61 491 -56
rect 512 -51 865 -31
rect 908 -36 960 -31
rect 512 -82 532 -51
rect 908 -56 918 -36
rect 938 -56 960 -36
rect 908 -59 960 -56
rect 260 -102 532 -82
<< via2 >>
rect 310 -5 330 15
rect 406 -4 426 16
rect 770 -10 790 10
<< metal3 >>
rect 401 16 441 21
rect 305 -5 310 15
rect 330 -5 353 15
rect 333 -36 353 -5
rect 401 -4 406 16
rect 426 -4 441 16
rect 401 -15 441 -4
rect 610 -10 770 10
rect 790 -10 795 10
rect 610 -36 630 -10
rect 333 -56 630 -36
<< labels >>
rlabel metal1 -45 77 -45 124 1 VDD!
rlabel metal1 -45 -124 -45 -77 1 VSS!
rlabel metal2 -24 -15 -24 15 1 C
rlabel metal3 401 -15 401 21 1 D
rlabel metal2 960 -59 960 -31 1 Q
rlabel metal1 101 -59 127 -33 1 nand1
rlabel metal1 223 59 249 59 1 nand0
rlabel metal2 496 36 496 62 1 nand3
rlabel metal1 666 28 666 59 1 nand2
rlabel metal1 881 59 911 59 1 nand5
rlabel metal1 66 -10 95 -10 1 R
<< end >>
